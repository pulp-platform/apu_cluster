`include "../ips/riscv/include/riscv_defines.sv"
