/scratch/gautschi/FP_PULP/pulp-dev/fe/rtl/includes/ulpsoc_defines.sv