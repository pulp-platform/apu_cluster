/scratch/gautschi/FP_PULP/pulp-dev/fe/ips/riscv/include/riscv_defines.sv