/scratch/gautschi/FP_PULP/pulp-dev/fe/rtl/includes/apu_defines.sv