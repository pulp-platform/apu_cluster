`ifdef SIMULATION
	`include "../ips/riscv/include/riscv_defines.sv"
`else 
	`include "riscv_defines.sv"
`endif
